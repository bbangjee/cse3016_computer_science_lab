`timescale 1ns / 1ps

module deMorganTwoB_tb;

reg a, b;
wire c;

deMorganTwoB test(
.a(a),
.b(b),

.c(c)
);

initial begin
  a = 1'b0;
  b = 1'b0;
  #160
  $finish;
end

always@(a or b) begin
  a <= #80 ~a;
  b <= #40 ~b;
end
    
endmodule
